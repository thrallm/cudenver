** Profile: "UniversalShiftReg-test_USR"  [ C:\Users\m\Desktop\CUDenver\github\cudenver\csci_1510\labs\lab06\final\lab06-final-pspicefiles\universalshiftreg\test_usr.sim ] 

** Creating circuit file "test_USR.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\Users\m\Desktop\CUDenver\github\cudenver\csci_1510\labs\lab06\final\lab06-final-pspicefiles\universalshiftreg\test_USR\tes"
+ "t_USR_profile.inc" 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\m\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 30ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\UniversalShiftReg.net" 


.END
