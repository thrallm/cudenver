** Profile: "test-D-from-JK-testDfromJK"  [ c:\users\m\desktop\cudenver\csci_1510\labs\lab05\lab05-pspicefiles\test-d-from-jk\testdfromjk.sim ] 

** Creating circuit file "testDfromJK.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../test-d-ff.stl" 
* From [PSPICE NETLIST] section of C:\Users\m\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\test-D-from-JK.net" 


.END
