** Profile: "half_adder_demo-halfadder"  [ C:\Users\m\Desktop\CUDenver\csci_1510\labs\lab04\lab04-PSpiceFiles\half_adder_demo\halfadder.sim ] 

** Creating circuit file "halfadder.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../xy.stl" 
.STMLIB "../../../2bitaddertest.stl" 
.STMLIB "../../../xy_carry_in.stl" 
* From [PSPICE NETLIST] section of C:\Users\m\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\half_adder_demo.net" 


.END
