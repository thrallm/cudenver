** Profile: "SCHEMATIC1-lab03_part1"  [ C:\Users\m\Desktop\CUDenver\csci_1510\labs\lab03\lab03-pspicefiles\schematic1\lab03_part1.sim ] 

** Creating circuit file "lab03_part1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../lab03_stimulus.stl" 
* From [PSPICE NETLIST] section of C:\Users\m\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
