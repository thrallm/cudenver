** Profile: "test_3bitReg-test_3bitparallelreg"  [ C:\Users\m\Desktop\CUDenver\github\cudenver\csci_1510\labs\lab06\parts\lab06-parts-pspicefiles\test_3bitreg\test_3bitparallelreg.sim ] 

** Creating circuit file "test_3bitparallelreg.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\Users\m\Desktop\CUDenver\github\cudenver\csci_1510\labs\lab06\parts\lab06-parts-pspicefiles\test_3bitreg\test_3bitparallel"
+ "reg\test_3bitparallelreg_profile.inc" 
* Local Libraries :
.STMLIB "C:/Users/m/Desktop/CUDenver/github/cudenver/csci_1510/labs/lab06/xyz.stl" 
* From [PSPICE NETLIST] section of C:\Users\m\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\test_3bitReg.net" 


.END
