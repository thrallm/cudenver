** Profile: "test_MUX-test_mux"  [ C:\Users\m\Desktop\CUDenver\github\cudenver\csci_1510\labs\lab06\parts\lab06-parts-pspicefiles\test_mux\test_mux.sim ] 

** Creating circuit file "test_mux.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
.INC "C:\Users\m\Desktop\CUDenver\github\cudenver\csci_1510\labs\lab06\parts\lab06-parts-pspicefiles\test_mux\test_mux\test_mux_pro"
+ "file.inc" 
* Local Libraries :
.STMLIB "C:/Users/m/Desktop/CUDenver/github/cudenver/csci_1510/labs/lab06/xyz.stl" 
* From [PSPICE NETLIST] section of C:\Users\m\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\test_MUX.net" 


.END
