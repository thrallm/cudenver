** Profile: "4to1MUX-xyz"  [ C:\USERS\THRALLM\DESKTOP\CSCI_1510\LABS\lab06\parts\lab06-parts-PSpiceFiles\4to1MUX\xyz.sim ] 

** Creating circuit file "xyz.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "C:/USERS/THRALLM/DESKTOP/CSCI_1510/LABS/lab06/xyz.stl" 
* From [PSPICE NETLIST] section of C:\Users\thrallm\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\4to1MUX.net" 


.END
